-----------------------------------------------------------------------
--  Robert Hana
--  CSUN Graduate Project ECE693, Spring 2019
--
--
--  File:               tb_AXISInjector.vhd
--  Description:        This file tests the AXI Sampler "TestSInjector_v1_0" 
--                      and is the basis IP for the AXI Sampler
----------------------------------------------------------------------------
--
--  Functional Tests Summary:
--      1. Test the AXI Reset in
--      2. SCRegister - Test R/W to the User registers 
--      3. SCRegister - Test Reset/Clear by User Register
--      4. SCRegister - Test enable/disable
--      5. SCRegister - Test Register gated sync-in (Injector has no gated sync-in)
--      6. Test non-gated sync-in                   (Deprecated feature.)
--      7. Test sticky flags (read when empty, write when full.)
--      8. Test single data writes.                 (Is tested by 7.)
--      9. Test Simple Burst writes                 (Is tested by 10.)
--      10.Test variety of burst write lengths from 4,8,16,32,64,128,256
----------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
  
--Work Dependencies
library work;
use work.axisampler_fifo_elegant_pkg.all; 
-- Uncomment the following library declaration if instantiating 
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity tb_AXIInjector is
--  Port ( ); Test bench as no ports!
end tb_AXIInjector;
 
architecture Behavioral of tb_AXIInjector is

 

            signal rd_clk                      :  std_logic                                                          := '0'           ;
            signal rd_clk_en                    : std_logic                                                          := '1'           ;
            signal dout                        :  std_logic_vector(31 downto 0)                                                       ;
            signal empty                        : std_logic                                                                           ;
            
            signal  rd_en                       :  std_logic                                                         := '0'           ;
          
                           -- Ports of Axi Slave Bus Interface S00_AXI_SamplerFIFO
                           
            signal s00_axi_samplerfifo_aclk    :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_aresetn :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_awid    :  std_logic_vector(C_S00_AXI_SamplerFIFO_ID_WIDTH-1 downto 0)       := "0"          ;
            signal s00_axi_samplerfifo_awaddr  :  std_logic_vector(C_S00_AXI_SamplerFIFO_ADDR_WIDTH-1 downto 0)     := "000000"     ;
            signal s00_axi_samplerfifo_awlen   :  std_logic_vector(7 downto 0)                                      := "00000000"   ;
            signal s00_axi_samplerfifo_awsize  :  std_logic_vector(2 downto 0)                                      := "000"        ;
            signal s00_axi_samplerfifo_awburst :  std_logic_vector(1 downto 0)                                      := "00"         ;
            signal s00_axi_samplerfifo_awlock  :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_awcache :  std_logic_vector(3 downto 0)                                      := "0000"       ;
            signal s00_axi_samplerfifo_awprot  :  std_logic_vector(2 downto 0)                                      := "000"        ;
            signal s00_axi_samplerfifo_awqos   :  std_logic_vector(3 downto 0)                                      := "0000"       ;
            signal s00_axi_samplerfifo_awregion:  std_logic_vector(3 downto 0)                                      := "0000"       ;
            signal s00_axi_samplerfifo_awuser  :  std_logic_vector(C_S00_AXI_SamplerFIFO_AWUSER_WIDTH-1 downto 0)                   ;
            signal s00_axi_samplerfifo_awvalid :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_awready :  std_logic                                                                         ;
            
            
            signal s00_axi_samplerfifo_wdata   :  std_logic_vector(C_S00_AXI_SamplerFIFO_DATA_WIDTH-1 downto 0)     := x"00000000"  ;
            signal s00_axi_samplerfifo_wstrb   :  std_logic_vector((C_S00_AXI_SamplerFIFO_DATA_WIDTH/8)-1 downto 0) := "0000"       ;
            signal s00_axi_samplerfifo_wlast   :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_wuser   :  std_logic_vector(C_S00_AXI_SamplerFIFO_WUSER_WIDTH-1 downto 0)                    ;
            signal s00_axi_samplerfifo_wvalid  :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_wready  :  std_logic                                                                         ;
            
            
            signal s00_axi_samplerfifo_bid     :  std_logic_vector(C_S00_AXI_SamplerFIFO_ID_WIDTH-1 downto 0)                       ;
            signal s00_axi_samplerfifo_bresp   :  std_logic_vector(1 downto 0)                                                      ;
            signal s00_axi_samplerfifo_buser   :  std_logic_vector(C_S00_AXI_SamplerFIFO_BUSER_WIDTH-1 downto 0)                    ;
            signal s00_axi_samplerfifo_bvalid  :  std_logic                                                                         ;
            signal s00_axi_samplerfifo_bready  :  std_logic                                                         := '0'          ;
            
            
            signal s00_axi_samplerfifo_arid    :  std_logic_vector(C_S00_AXI_SamplerFIFO_ID_WIDTH-1 downto 0)       := "0"          ;
            signal s00_axi_samplerfifo_araddr  :  std_logic_vector(C_S00_AXI_SamplerFIFO_ADDR_WIDTH-1 downto 0)     := "000000"     ;
            signal s00_axi_samplerfifo_arlen   :  std_logic_vector(7 downto 0)                                      := "00000000"   ;
            signal s00_axi_samplerfifo_arsize  :  std_logic_vector(2 downto 0)                                      := "000"        ;
            signal s00_axi_samplerfifo_arburst :  std_logic_vector(1 downto 0)                                      := "00"         ;
            signal s00_axi_samplerfifo_arlock  :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_arcache :  std_logic_vector(3 downto 0)                                      := "0000"       ;
            signal s00_axi_samplerfifo_arprot  :  std_logic_vector(2 downto 0)                                      := "000"        ;
            signal s00_axi_samplerfifo_arqos   :  std_logic_vector(3 downto 0)                                      := "0000"       ;
            signal s00_axi_samplerfifo_arregion    :  std_logic_vector(3 downto 0)                                  := "0000"       ;
            signal s00_axi_samplerfifo_aruser  :  std_logic_vector(C_S00_AXI_SamplerFIFO_ARUSER_WIDTH-1 downto 0)                   ;
            signal s00_axi_samplerfifo_arvalid :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_arready :  std_logic                                                                         ;
            
            
            signal s00_axi_samplerfifo_rid     :  std_logic_vector(C_S00_AXI_SamplerFIFO_ID_WIDTH-1 downto 0)       := "0"          ;
            signal s00_axi_samplerfifo_rdata   :  std_logic_vector(C_S00_AXI_SamplerFIFO_DATA_WIDTH-1 downto 0)                     ;  -- don't drive outputs in test bench
            signal s00_axi_samplerfifo_rresp   :  std_logic_vector(1 downto 0)                                      := "00"         ;
            signal s00_axi_samplerfifo_rlast   :  std_logic                                                         := '0'          ;    
            signal s00_axi_samplerfifo_ruser   :  std_logic_vector(C_S00_AXI_SamplerFIFO_RUSER_WIDTH-1 downto 0)                    ; 
            signal s00_axi_samplerfifo_rvalid  :  std_logic                                                         := '0'          ;
            signal s00_axi_samplerfifo_rready  :  std_logic                                                         := '0'          ;
      
     
            signal          sync_out            :  std_logic                                                                        ;
            --Test Bench Signals --
            
            type testBenchState is (test_none, test_axi_reset, test_user_regs, wait_for_interrupt,  test_enable_fifo, 
                                     test_write, test_fifo_reg_reset, test_fifo_internal_test, clearing_interrupt, test_enable, test_disable,
                                     test_enable_disable, test_correct_functioning, test_sticky_bits, test_burst_write, test_END);
                                     
            type testSubSection is (reset, enable, disable, idle, enable_and_reset, write, read, wait_for_interrupt, clearing_interrupt, write_burst);                                                             
            signal test : testBenchState := test_none;
            signal testSub : testSubSection := idle;
            signal EndOfTests : std_logic := '0';
            signal data : integer := 0;
            
            --an "Alias of a component, perhaps not supported by Xilinx.. --"
            --alias testVector is  uut.FIFOAXISlave_ins.fifo_inst.empty;
            --signal tvector : std_logic_vector(1 downto 0);
                   
begin

--------------------------------------------------------------------------------------
                           -- test bench clocks --
--------------------------------------------------------------------------------------                
        -- AXI Side Clock  --
        clocked_axi_process : process
        begin
            --200MHz AXI bus speed 2.5ns --
          wait for  2.5 ns; s00_axi_samplerfifo_aclk <= '0';
          wait for  2.5 ns; s00_axi_samplerfifo_aclk <= '1';
           data <= data + 1;
        end process;
        
        -- FIFO Sampler side Clock  -- 
        clocked_sampler_process: process
        begin
           --  ~83 MHz sampling speed 6ns per 1/2 period... or 12 ns period. (Some overflow possible still!)
            wait for 7 ns;  rd_clk <= '0';
            wait for 7 ns;  rd_clk <= '1';
           
        end process;

          uut : TestMultiReg_v1_0
          generic map(
            -- Users to add parameters here
            -- User parameters ends
            -- Do not modify the parameters beyond this line
            -- Parameters of AXI4 Slave Bus Interface S00_AXI
            -- Parameters of Axi Slave Bus Interface S00_AXI_SamplerFIFO
            C_S00_AXI_ID_WIDTH      =>   C_S00_AXI_SamplerFIFO_ID_WIDTH ,
            C_S00_AXI_DATA_WIDTH    =>   C_S00_AXI_SamplerFIFO_DATA_WIDTH,
            C_S00_AXI_ADDR_WIDTH    =>   C_S00_AXI_SamplerFIFO_ADDR_WIDTH,
            C_S00_AXI_AWUSER_WIDTH  =>   C_S00_AXI_SamplerFIFO_AWUSER_WIDTH,
            C_S00_AXI_ARUSER_WIDTH  =>   C_S00_AXI_SamplerFIFO_ARUSER_WIDTH,
            C_S00_AXI_WUSER_WIDTH   =>   C_S00_AXI_SamplerFIFO_WUSER_WIDTH,
            C_S00_AXI_RUSER_WIDTH   =>   C_S00_AXI_SamplerFIFO_RUSER_WIDTH,
            C_S00_AXI_BUSER_WIDTH   =>   C_S00_AXI_SamplerFIFO_BUSER_WIDTH

          )
          port map(

		    -- Users to add ports here
           -- FIFO signals --
          
           trigger_out                  =>              sync_out                   ,
           rd_clk                       =>              rd_clk                     ,
           rd_clk_en                    =>              rd_clk_en                  , 
           dout                         =>              dout                       , 
           empty                        =>              empty                      ,    
            -- User ports ends
            -- Do not modify the ports beyond this line
            s00_axi_aclk    =>              s00_axi_samplerfifo_aclk    ,
            s00_axi_aresetn =>              s00_axi_samplerfifo_aresetn ,
            s00_axi_awid    =>              s00_axi_samplerfifo_awid    ,
            s00_axi_awaddr  =>              s00_axi_samplerfifo_awaddr  ,
            s00_axi_awlen   =>              s00_axi_samplerfifo_awlen   ,
            s00_axi_awsize  =>              s00_axi_samplerfifo_awsize  ,
            s00_axi_awburst =>              s00_axi_samplerfifo_awburst ,
            s00_axi_awlock  =>              s00_axi_samplerfifo_awlock  ,
            s00_axi_awcache =>              s00_axi_samplerfifo_awcache ,
            s00_axi_awprot  =>              s00_axi_samplerfifo_awprot  ,
            s00_axi_awqos   =>              s00_axi_samplerfifo_awqos   ,
            s00_axi_awregion    =>          s00_axi_samplerfifo_awregion    ,
            s00_axi_awuser  =>              s00_axi_samplerfifo_awuser  ,
            s00_axi_awvalid =>              s00_axi_samplerfifo_awvalid ,
            s00_axi_awready =>              s00_axi_samplerfifo_awready ,
            s00_axi_wdata   =>              s00_axi_samplerfifo_wdata   ,
            s00_axi_wstrb   =>              s00_axi_samplerfifo_wstrb   ,
            s00_axi_wlast   =>              s00_axi_samplerfifo_wlast   ,
            s00_axi_wuser   =>              s00_axi_samplerfifo_wuser   ,
            s00_axi_wvalid  =>              s00_axi_samplerfifo_wvalid  ,
            s00_axi_wready  =>              s00_axi_samplerfifo_wready  ,
            s00_axi_bid     =>              s00_axi_samplerfifo_bid ,
            s00_axi_bresp   =>              s00_axi_samplerfifo_bresp   ,
            s00_axi_buser   =>              s00_axi_samplerfifo_buser   ,
            s00_axi_bvalid  =>              s00_axi_samplerfifo_bvalid  ,
            s00_axi_bready  =>              s00_axi_samplerfifo_bready  ,
            s00_axi_arid    =>              s00_axi_samplerfifo_arid    ,
            s00_axi_araddr  =>              s00_axi_samplerfifo_araddr  ,
            s00_axi_arlen   =>              s00_axi_samplerfifo_arlen   ,
            s00_axi_arsize  =>              s00_axi_samplerfifo_arsize  ,
            s00_axi_arburst =>              s00_axi_samplerfifo_arburst ,
            s00_axi_arlock  =>              s00_axi_samplerfifo_arlock  ,
            s00_axi_arcache =>              s00_axi_samplerfifo_arcache ,
            s00_axi_arprot  =>              s00_axi_samplerfifo_arprot  ,
            s00_axi_arqos   =>              s00_axi_samplerfifo_arqos   , 
            s00_axi_arregion    =>          s00_axi_samplerfifo_arregion,
            s00_axi_aruser  =>              s00_axi_samplerfifo_aruser  ,
            s00_axi_arvalid =>              s00_axi_samplerfifo_arvalid ,
            s00_axi_arready =>              s00_axi_samplerfifo_arready ,
            
            
            s00_axi_rid     =>              s00_axi_samplerfifo_rid     ,
            s00_axi_rdata   =>              s00_axi_samplerfifo_rdata   ,
            s00_axi_rresp   =>              s00_axi_samplerfifo_rresp   ,
            s00_axi_rlast   =>              s00_axi_samplerfifo_rlast   ,
            s00_axi_ruser   =>              s00_axi_samplerfifo_ruser   ,
            s00_axi_rvalid  =>              s00_axi_samplerfifo_rvalid  ,
            s00_axi_rready  =>              s00_axi_samplerfifo_rready  

        
          );        
        
    --procedures can drive signals if they are in a process without a sensitivity list
    -- This is how the code should be ordered!
    -- we can have more than one process like this!!! So it can handle different signals concurrently

    -- This is the overall Test Process here --
    test_this : process
    
        variable  writes       : integer := 0  ;
        variable  waitClocks   : integer := 0  ;
        variable  writeRegAddr : integer := 0  ;
        variable  readRegAddr  : integer := 0  ;
        variable  dataValue    : integer := 123;
       
        variable resetCount    : integer := 0;
        
    
    begin    
    
        --------------------------------- No test  ------------------------------
        -- Start without a test and without reset asserted
        -- There should be a few unknown signals going on here.
        test <= test_none;
        testSub <= idle;
        s00_axi_samplerfifo_aresetn <= '1'; 
        waitClocks := 100; 
        wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
        

        --------------------------------- 1. Test AXI Reset ------------------------------
        -- Notes: testing whether or not the axi global reset will reset the device
        test <= test_axi_reset; 
        testSub <= idle;
        s00_axi_samplerfifo_aresetn <= '1';
        waitClocks := 50;  
        wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
        
        testSub <= reset;
        resetCount := 0;
        for i in 0 to 16 loop
            s00_axi_samplerfifo_aresetn <= '0';
            wait until rising_edge(s00_axi_samplerfifo_aclk);
            resetCount := resetCount  + 1;
        end loop;
        report "Reset is asserted for " & integer'image(resetCount) & " clock cycles." severity note;
        assert (resetCount >= 16 ) report "AXI Global Reset must be asserted at least an N = 16 number of write clock cycles or read clocks of the slowest clock, generally for Xilinx IP" severity failure;
           
        test <= test_none;
        testSub <= idle;
        s00_axi_samplerfifo_aresetn <= '1'; 
        waitClocks := 25; 
        wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
        
       ------------------- End Test AXI Reset ----------------------------------------

      
        
             
        ---------------------------------   2. Test SCRegister - Test R/W to the User registers ------------------------
        -- verify writing can be done to the other 3 registers (without enabling or disabling. So don't touch the upper 6 bits)
        -- <128,192>, <256,384>, <384,576>
        -- Verify sync_out goes high when read_enable is high.
          test <= test_user_regs;
          testSub <= idle;
          for i in 1 to 3 loop
              waitClocks := 75; 
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
             --do something else if write isn't enabled, ...lets read and write to the AXISlave registers.
              waitClocks := 10; 
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
             

              -- Write data to the registers --
              testSub <= write;
              dataValue    := 128 * i;
              writeRegAddr := 4  ;
              write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                  s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                  s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
                                 
              dataValue    := 192 * i;
              writeRegAddr := 8  ;
              write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                  s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                  s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
                
              -- Then read the data back out --
              testSub <= read;
              waitClocks := 50; 
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
             
              readRegAddr := 4;
              read_from_register(readRegAddr,  s00_axi_samplerfifo_aclk , s00_axi_samplerfifo_araddr, s00_axi_samplerfifo_arvalid , s00_axi_samplerfifo_arlen ,s00_axi_samplerfifo_arsize , s00_axi_samplerfifo_rready );
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
             
              readRegAddr := 8;
              read_from_register(readRegAddr,  s00_axi_samplerfifo_aclk , s00_axi_samplerfifo_araddr, s00_axi_samplerfifo_arvalid , s00_axi_samplerfifo_arlen ,s00_axi_samplerfifo_arsize , s00_axi_samplerfifo_rready );
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
         
              waitClocks := 50; 
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
    
          end loop;
          
          ---------------------------------   END  Test SCRegister - Test R/W to the User registers ------------------------
    
            
            
            --------------------------------- 3. SCRegister - Test Reset/Clear by User Register------------------------  
            -- Notes: Tests writing to the SCRegister all lower 6 bits and verify they clear
            
            
          test <= test_user_regs;
          testSub <= idle;
            for i in 1 to 3 loop
                waitClocks := 75; 
                wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
               --do something else if write isn't enabled, ...lets read and write to the AXISlave registers.
                waitClocks := 10; 
                wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
               
  
                -- Write data to the registers --
                testSub <= write;
                dataValue    := 127;
                writeRegAddr := 4  ;
                write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                    s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                    s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
  
                -- Then read the data back out --
                waitClocks := 50; 
                wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
               testSub <= read;
                readRegAddr := 4;
                read_from_register(readRegAddr,  s00_axi_samplerfifo_aclk , s00_axi_samplerfifo_araddr, s00_axi_samplerfifo_arvalid , s00_axi_samplerfifo_arlen ,s00_axi_samplerfifo_arsize , s00_axi_samplerfifo_rready );
                wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);

                testSub <= idle;
                waitClocks := 250; 
                wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
                
                testSub <= read;
                readRegAddr := 4;
                read_from_register(readRegAddr,  s00_axi_samplerfifo_aclk , s00_axi_samplerfifo_araddr, s00_axi_samplerfifo_arvalid , s00_axi_samplerfifo_arlen ,s00_axi_samplerfifo_arsize , s00_axi_samplerfifo_rready );
                wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);

           
                waitClocks := 50; 
                wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
      
            end loop;
            
             --------------------------------- END  SCRegister - Test Reset/Clear by User Register------------------------ 

            
            
            --------------------------------- 4. Test SCRegister - Test enable/disable  ---------------------------------
            --  Notes: The AXI fifo is loaded with data. 
            --         The enable/disable is tested. When enabled, data should be read out
            --          When disabled, data won't be read out. Data not read out hangs on the data output.
            
             test <= test_enable_disable;
             testSub <= idle;
              waitClocks := 10; 
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
              --write some data to it
              testSub <= write;
              for i in 1 to 100 loop
                  dataValue    := i ;
                  writeRegAddr := 0  ;
                  write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                      s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                      s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
              end loop;
              
              testSub <= idle;
              waitClocks := 10; 
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
              
              for i in 1 to 5 loop
              
                  test <= test_enable;
                  --enable it--
                  testSub <= enable;
                  dataValue    := 2 ;
                  writeRegAddr := 4  ;
                  write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                      s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                      s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
                  waitClocks := 100; 
                  wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);                                 
                                      
                  test <= test_disable;  
                  testSub <= disable;                
                  --disable it--
                  dataValue    := 0 ;
                  writeRegAddr := 4 ;
                  write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                      s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                      s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        ); 
                  waitClocks := 100; 
                  wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);                                      
              end loop;

              ---------------------------- END Test SCRegister - Test enable/disable -------------------------------------------------------
              
              
              --      5. SCRegister - Test Register gated sync-in (Injector has no gated sync-in) No Test.
              --      6. Test non-gated sync-in                                                   (Deprecated feature.)
              
              --------------------------            7. Test sticky flags (read when empty, write when full.) -------------------------------
              -- Notes: Sticky bits return 0x6 when overflow ocurred and enabled, returns 12 after disabled 0xC 
               test <= test_sticky_bits;  
               testSub <= idle; 
               waitClocks := 10; 
               wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
               
               --reset it
               testSub <= reset;
               dataValue    := 1;
               writeRegAddr := 4  ;
               write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                   s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                   s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
               waitClocks := 300;                 
               wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);  
               
               
               -- read SC register
               testSub <= read;
               readRegAddr := 4;
               read_from_register(readRegAddr,  s00_axi_samplerfifo_aclk , s00_axi_samplerfifo_araddr, s00_axi_samplerfifo_arvalid , s00_axi_samplerfifo_arlen ,s00_axi_samplerfifo_arsize , s00_axi_samplerfifo_rready );
               wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
               
               
               --enable before writing data to it
               testSub <= enable;
               dataValue    := 2;
               writeRegAddr := 4  ;
               write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                   s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                   s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
               
               
               --wait for some time..this should cause Underflow flag to go high.
               waitClocks := 300;                 
               wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk); 
               
               --read sc register
               testSub <= read;
               readRegAddr := 4;
               read_from_register(readRegAddr,  s00_axi_samplerfifo_aclk , s00_axi_samplerfifo_araddr, s00_axi_samplerfifo_arvalid , s00_axi_samplerfifo_arlen ,s00_axi_samplerfifo_arsize , s00_axi_samplerfifo_rready );
               wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
               
               
               
               --disable it before writing data to it
               testSub <= enable;
               dataValue    := 0;
               writeRegAddr := 4  ;
               write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                   s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                   s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
                                   
               --write too much to it
               for i in 0 to 2200 loop
                   dataValue    := i;
                   writeRegAddr := 0  ;
                   write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                       s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                       s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
               
               end loop;
               
               
               
               --read sc register
               readRegAddr := 4;
               read_from_register(readRegAddr,  s00_axi_samplerfifo_aclk , s00_axi_samplerfifo_araddr, s00_axi_samplerfifo_arvalid , s00_axi_samplerfifo_arlen ,s00_axi_samplerfifo_arsize , s00_axi_samplerfifo_rready );
               wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
               
               
               --reset it
                 testSub <= reset;
                 dataValue    := 1;
                 writeRegAddr := 4  ;
                 write_to_register(  dataValue, writeRegAddr,  s00_axi_samplerfifo_aclk                                                                                                  , 
                                     s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                                     s00_axi_samplerfifo_wdata ,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
                 waitClocks := 300;                 
                 wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);                    
               --read sc register
               
               ----------------------------  End Test sticky flags (read when empty, write when full.)-------------------------------------------------------
              
              
              -------------                 9. and 10.  Test  Burst writes     ----------------------
               test <= test_burst_write;  
               for i in 2 to 8 loop
                 testSub <= write_burst; 
                 writeRegAddr := 0  ;
                 writes := 2**i;
                 write_axi_slave(   writeRegAddr, data, writes,  s00_axi_samplerfifo_aclk                                                                             , 
                          s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                           s00_axi_samplerfifo_wdata, s00_axi_samplerfifo_wready,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
                           
                 testSub <= idle;          
                 waitClocks := 300;                 
                 wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
                end loop ;
              
             ----- Last bursts
             testSub <= write_burst; 
             writeRegAddr := 0  ;
             for i in 1 to 4 loop
             writes := 4;
             write_axi_slave(   writeRegAddr, data, writes,  s00_axi_samplerfifo_aclk                                                                             , 
                      s00_axi_samplerfifo_awaddr, s00_axi_samplerfifo_awvalid,  s00_axi_samplerfifo_awlen  , s00_axi_samplerfifo_awsize                                   ,  
                       s00_axi_samplerfifo_wdata, s00_axi_samplerfifo_wready,  s00_axi_samplerfifo_wvalid,  s00_axi_samplerfifo_wlast , s00_axi_samplerfifo_wstrb,  s00_axi_samplerfifo_bready        );
                   
              end loop;
              
              
              test <= test_END;
              EndOfTests <= '1';
              testSub <= idle;

              assert false report "writes value on burst length are always (writes + 1.) so if length is 0, then 1 read is implied." severity note;
              assert false report "Reset must be asserted for an N = 16 number of write clock cycles or read clocks, here its done with a counter internally for the register reset." severity note;
              assert false report "writes value on burst length are always (writes + 1.) so if length is 0, then 1 read is implied." severity note;
              assert false report "Reset must be asserted for an N = 16 number of write clock cycles or read clocks, here its done with a counter internally for the register reset." severity note;   
              waitClocks := 100; 
              wait_for_clock_cycles(waitClocks,s00_axi_samplerfifo_aclk);
              wait;


            --Conclusion: If you enable it and then start writing to it (instead of writing to it first, and then enabling it), the data coming out will not occor on
            -- every read cycle because it may take a couple of the write_clock cycles to get the data IN, and the read/write pointers in the FIFO are going to be
            --right on top of each other... this will happen read/write clocks that are close in frequency and bursts are not used, and this can be a problem. The device should first
            --be reset.. next written to... next enabled... .. and then the Zynq processor should wait for the interrupt before providing a burst write. Without
            -- doing these things in this order... there could be data corruption (essentially trying to read from it while it is empty.)
            
            -- Read the Data from the Fifo -- (should be able to handle 256 words per burst.)
            
            --Contiguous writes working fine for multiple burst writes up to 2047, 
            --                .. size 2048 or higher results in reading from an empty fifo, with junk data x"00000000" in simulation
            --   The read/write flag status should be verified in hardware
            --   It is reasonable there is a 1 clock cycle delay before empty flag is asserted.
            --   It doesn't make sense the depth is 2047 and not 2048 (so this is an issue that needs to be explored.)
            --FIFO Size is 2048, when writes = 0, writes 1 time... read size is actually ""writes + 1"  128 x 15 = 1920 ; "127" is actually "128" because if it was "0" it would be "1" ..so add 1.

           
    

    end process;

    
    ---   
    



end Behavioral;


